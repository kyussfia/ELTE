6
1
000000
000200
001000
002000
000000
000000
000
00000000000000
00000000000000
00000000000000
00000002000000
00000000000000
00000010000000
00000000000000
00000000000000
00000000000000
00000000000000
00000000000000
